`timescale 1ns / 1ps

module comp_fp4(
    input logic [3:0] E1,E2,E3,C,
    input logic [3:0] d41,d42,d51,d52,d61,d62,           //connect 6th block in top module
    output logic [3:0] Emax
    );
    
   // no need pf this module
    
endmodule
